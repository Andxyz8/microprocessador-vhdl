LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY rom IS
    PORT
    (
        clk     : IN STD_LOGIC;
        read    : IN STD_LOGIC;
        address : IN UNSIGNED (6 DOWNTO 0); -- Verificar a quantidade exata depois
        data    : OUT UNSIGNED (14 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE a_rom OF rom IS
    TYPE mem IS ARRAY (0 TO 127) OF UNSIGNED(14 DOWNTO 0);
    CONSTANT conteudo_rom : mem := (                            --  
        0       => B"110000_001_000111",     -- LD $R1, 7       --  0 + 7   1 0
        1       => B"001000_001_000111",     -- LD (0x7), $R1   --  0 + r1  0 0
        2       => B"011000_010_000111",     -- LD $R2, (0x7)   --  0x + 0  0 1
        3       => B"000000_000_000000",     --
        4       => B"000000_000_000000",     --
        5       => B"000000_000_000000",     --
        6       => B"000000_000_000000",     --
        15      => B"000000_000_000000",     --
        OTHERS  => (OTHERS => '0')
    );
    
BEGIN
    PROCESS(clk)
    BEGIN
        IF (read = '1') THEN
            IF(rising_edge(clk)) THEN
                data <= conteudo_rom(TO_INTEGER(address));
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE a_rom;
